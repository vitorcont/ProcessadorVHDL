LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY mem IS
PORT(
	address: in integer range 0 to 8;
	data: out STD_LOGIC_VECTOR(17 downto 0));
END mem;

ARCHITECTURE Behavior OF mem IS
	type memoria is array (0 to 8) of STD_LOGIC_VECTOR (17 downto 0);
	constant rom: memoria := ( 
	"100000100000001000", "100100000000101000", "101000000000010001", "001101000000000001", 
	"010000000100000100", "010110001100000011", "011000100000000010", "011101110000000100", "000000000000000000"
	);
	BEGIN
		data <= rom(address);
END Behavior;