LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RegInst IS
PORT(
	Instruction : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	Op 		: OUT STD_LOGIC ;
	FUNC	: OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
	AdressA 	:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
	AdressB 	:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
	WriteAdress 	:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
	IMED 	:	OUT	STD_LOGIC_VECTOR(7 DOWNTO 0);
	Clock 	: IN STD_LOGIC );
END RegInst;

ARCHITECTURE Behavior OF RegInst IS
	SIGNAL R1	:	STD_LOGIC_VECTOR(17 DOWNTO 0);
	-- Alterar do Clock
	BEGIN
			R1<=Instruction;
			Op <=R1(17);
			FUNC<=R1(2 DOWNTO 0);
			AdressA<=R1(13 DOWNTO 11);
			AdressB<=R1(10 DOWNTO 8);
			WriteAdress<=R1(16 DOWNTO 14);
			IMED<=R1(10 DOWNTO 3);
END Behavior;