LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MUX IS
PORT(
	Banco	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	Imed	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	IMEDSrc 	: IN STD_LOGIC;
	FinalValue 	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END MUX;

ARCHITECTURE Behavior OF MUX IS
BEGIN
	PROCESS(IMEDSrc,Banco,Imed)
		BEGIN
			IF IMEDSrc = '0' THEN
				FinalValue <= Banco;
			ELSE
				FinalValue <= Imed;
			END IF;
	END PROCESS;
END Behavior;